$display("NPU init done.");
$display("Weight loaded.");
$display("Input loaded.");
h2f_pio32=32'hc0000000;h2f_write=1;@(negedge clk)h2f_write=0;
@(posedge |(f2h_pio32 & 32'h10000000));@(negedge clk);
$display("Fetch done.");
h2f_pio32=32'ha6;h2f_write=1;@(negedge clk)h2f_write=0;
@(posedge |(f2h_pio32 & 32'h40000000));@(negedge clk);
$display("Load done.");
h2f_pio32=32'h80080001;h2f_write=1;@(negedge clk)h2f_write=0;
@(posedge |(f2h_pio32 & 32'h80000000));@(negedge clk);
$display("Move done.");
h2f_pio32=32'he0000000;h2f_write=1;@(negedge clk)h2f_write=0;
@(posedge |(f2h_pio32 & 32'h1));@(negedge clk);
$display("Exec done.");
h2f_pio32=32'ha0829c01;h2f_write=1;@(negedge clk)h2f_write=0;
@(posedge |(f2h_pio32 & 32'h80000000));@(negedge clk);
$display("Move done.");
h2f_pio32=32'h54f00001;h2f_write=1;@(negedge clk)h2f_write=0;
@(posedge |(f2h_pio32 & 32'h40000000));@(negedge clk);
$display("Store done.");
